module mux8to1 (
    input  [7:0] d,
    input  [2:0] sel,
    output reg y          
);
    always @(*) begin
        case (sel)
            3'b000: y = d[0];
            3'b001: y = d[1];
            3'b010: y = d[2];
            3'b011: y = d[3];
            3'b100: y = d[4];
            3'b101: y = d[5];
            3'b110: y = d[6];
            3'b111: y = d[7];
            default: y = 1'b0;
        endcase
    end
endmodule

`timescale 1ns/1ps
module tb_mux8to1;
    reg  [7:0] d;     
    reg  [2:0] sel;    
    wire y;            
    mux8to1 uut (
        .d(d),
        .sel(sel),
        .y(y)
    );

    integer i;
    initial begin
        $display("Sel\tD\t\tY");
        $monitor("%b\t%b\t%b", sel, d, y);

        // Test 16 cases: each input bit once with 0, once with 1
        for (i = 0; i < 8; i = i + 1) begin
            sel = i;              // Select input i
            
            // Case 1: input bit = 0
            d = 8'b0;             // all 0s
            #5;

            // Case 2: input bit = 1
            d = (1 << i);         // only d[i] = 1
            #5;
        end

        #10 $finish;
    end
    initial begin
        $dumpfile("mux.vcd");
        $dumpvars(0,tb_mux8to1);
    end
endmodule