module not_from_nor(
    input a,
    output y
    );
    nor (y, a, a);
endmodule